library ieee;
 use ieee.std_logic_1164.all;
 use ieee.std_logic_misc.all;
 use ieee.numeric_std.all;
 use work.Constants.all;
 use work.Types.all;
 package Arrays0_0000 is
 constant initPredict : ty := to_ty(0);
 constant feature : intArray(nNodes-1 downto 0)  :=  (1,72,72,10,7,405,122,377,377,81,81,5,72,377,22,404,404,221,7,404,7,85,19,22,395,10,22,404,404,14,8,42,363,-2,407,139,120,424,446,22,384,29,373,1,7,19,81,54,404,-2,81,-2,5,22,81,147,404,7,22,-2,-2,54,72,471,-2,377,-2,-2,-2,424,81,64,93,377,-2,332,395,439,396,81,395,7,-2,424,43,64,-2,-2,182,144,404,43,395,377,388,371,-2,346,396,43,43,368,54,395,402,396,143,417,404,1,143,377,402,-2,-2,-2,3,-2,-2,0,368,388,404,147,-2,-2,86,-2,-2,391,404,95,-2,363,-2,59,64,-2,-2,-2,-2,148,149,8,402,395,373,20,-2,319,402,90,373,7,439,42,215,321,-2,404,-2,-2,-2,20,416,215,8,411,42,65,111,-2,-2,-2,-2,93,165,-2,122,416,402,-2,120,294,8,321,-2,-2,-2,368,42,321,365,-2,8,384,5,-2,-2,404,439,23,321,381,3,391,-2,-2,313,313,-2,139,-2,19,72,-2,313,144,108,402,-2,233,164,232,214,446,388,-2,72,-2,-2,402,120,-2,-2,-2,465,391,214,360,62,-2,-2,-2,65,-2,-2,405,407,-2,-2,57,327,144,27,321,72,-2,-2,-2,364,424,364,72,72,-2,-2,-2,22,27,315,471,364,214,363,411,313,391,72,-2,72,19,471,19,72,0,19,7,396,-2,-2,-2,-2,315,-2,407,72,-2,-2,-2,384,396,411,144,391,402,-2,-2,-2,417,397,14,-2,-2,149,-2,-2,23,-2,364,377,391,214,-2,-2,8,-2,-2,-2,396,-2,143,214,72,365,-2,-2,-2,-2,-2,-2,-2,-2,315,-2,-2,-2,22,143,72,-2,396,353,439,454,93,-2,-2,-2,396,402,365,214,63,-2,-2,365,72,360,-2,-2,-2,-2,402,-2,143,-2,-2,-2,-2,-2,65,347,441,-2,-2,-2,-2,-2,377,-2,-2,-2,-2,313,446,20,364,411,-2,377,363,-2,-2,-2,377,-2,-2,-2,-2,-2,-2,-2,14,10,365,365,377,-2,149,353,165,93,-2,-2,346,394,-2,417,-2,144,-2,-2,391,-2,313,8,377,-2,231,-2,377,-2,143,143,11,-2,-2,-2,377,-2,-2,-2,-2,-2,-2,-2,397,-2,-2,388,-2,371,-2,139,-2,72,-2,-2,-2,-2,7,-2,64,364,19,-2,64,368,1,-2,-2,-2,294,397,-2,-2,-2,-2,-2,-2,45,215,-2,7,-2,-2,63,395,-2,395,-2,-2,-2,424,-2,-2,-2,0,397,-2,407,395,182,122,388,-2,360,14,364,395,381,14,364,-2,7,-2,138,-2,-2,319,1,-2,-2,395,-2,-2,-2,353,27,22,5,395,-2,-2,72,388,165,65,-2,377,-2,397,-2,-2,-2,0,7,360,-2,-2,5,43,0,62,396,381,-2,404,45,1,424,-2,-2,-2,-2,381,377,-2,377,-2,-2,-2,-2,-2,86,3,313,90,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2,-2);
 constant threshold_int : intArray(nNodes-1 downto 0)  :=  (-14360,-4083,-13993,11903,512,-10240,213,11327,-15694,-8751,11785,-1655,9827,-7756,11700,-12275,-1272,3605,-1844,0,15107,3511,-1182,-15843,-8332,-4171,209,1119,-9504,11777,-1999,-12635,-2552,0,6144,-9449,-11905,-541,3584,-14247,-4608,-10991,512,-11500,-4628,-13945,-1896,-809,15360,0,-8372,0,-96,7786,-10761,-9887,10487,5873,13689,0,0,953,-10560,512,0,11788,0,0,0,-8435,1160,1814,3263,-11098,0,9490,-8936,-10240,5120,-5667,6594,10255,0,-5990,0,-11444,0,0,11464,-5768,-3606,-8710,3818,11920,-15014,512,0,-4348,9000,3584,5667,-10649,0,10485,14405,5555,-7914,-11059,15790,920,-8099,3460,752,0,0,0,-11235,0,0,-15796,-13917,-1039,15360,1536,0,0,96,0,0,787,11910,6505,0,-7825,0,14179,7962,0,0,0,0,13132,11689,14019,-9216,10326,512,7279,0,-7061,6817,5986,512,-7806,7168,-225,15064,-12899,0,11422,0,0,0,7647,9728,-8490,-15082,-11262,-1199,-1473,-13823,0,0,0,0,-12114,-11320,0,-14307,4067,-12288,0,-8866,12662,2839,-4468,0,0,0,2734,7159,-1971,14848,0,-11553,-4048,-9806,0,0,-12833,3584,8704,358,-4503,7153,-5090,0,0,-4896,6891,0,11947,0,5671,7177,0,10949,10214,3362,-10014,0,7719,6649,9216,-7989,3584,-9541,0,6646,0,0,512,-9041,0,0,0,512,13460,-11405,-9124,10241,0,0,0,4880,0,0,-2048,-14336,0,0,2592,-12629,6712,5565,9956,-4493,0,0,0,12641,1371,-9728,12011,7879,0,0,0,7962,-4373,12228,512,-6572,8723,-6656,15129,512,-3026,571,0,8315,-14884,512,9381,-8870,-2798,2707,4765,-4081,0,0,0,0,-15718,0,-5940,12467,0,0,0,4969,9749,11497,10602,-14695,-5671,0,0,0,6656,1996,4599,0,0,1212,0,0,-7391,0,3822,571,7911,13638,0,0,13569,0,0,0,4054,0,-301,-2771,8333,3031,0,0,0,0,0,0,0,0,1766,0,0,0,11328,2316,-8582,0,797,-494,4096,512,3153,0,0,0,-5175,2591,10064,-5043,8357,0,0,9883,-2288,-4315,0,0,0,0,4954,0,15195,0,0,0,0,0,-7596,-1400,4608,0,0,0,0,0,-12695,0,0,0,0,14715,-4096,-1128,-13242,13312,0,-2270,-6313,0,0,0,4743,0,0,0,0,0,0,0,-1004,2048,-7622,-513,8135,0,15519,7943,3358,-6584,0,0,-7134,14593,0,-11264,0,-8990,0,0,11477,0,-11902,4549,-12632,0,1833,0,-6183,0,6921,-10401,30,0,0,0,-2250,0,0,0,0,0,0,0,-7553,0,0,7540,0,512,0,-13421,0,8083,0,0,0,0,-5229,0,-1777,2426,-5755,0,-7550,-12300,-14462,0,0,0,9165,10272,0,0,0,0,0,0,-40,-3885,0,-5804,0,0,708,-2482,0,5933,0,0,0,730,0,0,0,-3950,11836,0,-6656,-5936,-10159,-9510,12595,0,-6137,4683,-3367,5162,13090,12328,3500,0,-6086,0,-12560,0,0,-210,9285,0,0,15754,0,0,0,10559,2340,4131,4548,1793,0,0,-2030,7734,1222,-3059,0,10646,0,-15004,0,0,0,196,7937,-13238,0,0,8002,6567,-11282,13336,4485,13939,0,6296,13241,-3548,0,0,0,0,0,12351,12064,0,-8382,0,0,0,0,0,-2177,-6221,-9233,9742,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024,-1024);
 constant children_left : intArray(nNodes-1 downto 0)  :=  (1,3,5,7,11,9,13,15,27,17,29,25,21,19,23,31,59,33,61,57,53,35,55,51,49,47,45,43,39,37,41,63,113,733,65,115,111,107,67,109,105,103,101,99,97,93,69,95,91,735,89,737,87,85,83,81,79,77,75,739,741,73,71,117,743,197,745,747,749,119,199,195,191,121,751,193,189,187,185,183,181,177,753,123,179,175,755,757,173,171,169,167,165,163,161,159,759,157,155,153,151,147,125,149,145,143,141,139,137,135,133,131,129,761,763,765,127,767,769,201,307,203,309,305,771,773,301,775,777,205,303,299,779,297,781,295,293,783,785,787,789,291,287,207,289,285,283,281,791,279,277,275,273,271,269,267,265,263,793,261,795,797,799,257,209,259,255,253,251,249,247,801,803,805,807,245,243,809,241,239,237,811,235,233,231,229,813,815,817,227,225,223,221,819,219,217,215,821,823,213,211,311,453,313,455,451,825,827,447,315,829,449,831,445,443,833,441,439,437,433,835,317,435,431,429,427,425,837,423,839,841,421,419,843,845,847,417,415,413,411,409,849,851,853,407,855,857,403,319,859,861,405,401,399,397,395,393,863,865,867,391,389,387,385,383,869,871,873,381,379,377,375,373,371,369,367,365,363,361,875,359,357,355,353,351,349,347,345,341,877,879,881,883,321,885,343,339,887,889,891,337,335,333,331,329,327,893,895,897,325,323,457,899,901,587,903,905,459,907,589,585,581,461,909,911,583,913,915,917,579,919,577,575,573,571,921,923,925,927,929,931,933,935,567,937,939,941,463,569,565,943,563,561,559,557,555,945,947,949,553,551,549,547,545,951,953,543,541,537,955,957,959,961,465,963,539,965,967,969,971,973,535,533,531,975,977,979,981,983,529,985,987,989,991,527,525,523,521,519,993,517,515,995,997,999,513,1001,1003,1005,1007,1009,1011,1013,511,509,507,505,503,1015,501,499,497,495,1017,1019,493,491,1021,489,1023,487,1025,1027,485,1029,483,481,479,1031,475,1033,467,1035,477,473,471,1037,1039,1041,469,1043,1045,1047,1049,1051,1053,1055,591,1057,1059,729,1061,593,1063,731,1065,727,1067,1069,1071,1073,723,1075,595,725,721,1077,719,717,715,1079,1081,1083,713,709,1085,1087,1089,1091,1093,1095,597,711,1097,707,1099,1101,705,703,1103,701,1105,1107,1109,699,1111,1113,1115,697,695,1117,693,691,689,687,685,1119,683,679,599,681,677,675,673,1121,671,1123,669,1125,1127,667,665,1129,1131,663,1133,1135,1137,661,659,657,655,653,1139,1141,651,649,647,645,1143,643,1145,641,1147,1149,1151,639,637,635,1153,1155,633,631,629,627,625,623,1157,621,617,601,619,1159,1161,1163,1165,615,613,1167,611,1169,1171,1173,1175,1177,609,607,605,603,1179,1181,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,1183,1185,1187,1189,1191,1193,1195,1197,1199,1201,1203,1205,1207,1209,1211,1213,1215,1217,1219,1221,1223,1225,1227,1229,1231,1233,1235,1237,1239,1241,1243,1245,1247,1249,1251,1253,1255,1257,1259,1261,1263,1265,1267,1269,1271,1273,1275,1277,1279,1281,1283,1285,1287,1289,1291,1293,1295,1297,1299,1301,1303,1305,1307,1309,1311,1313,1315,1317,1319,1321,1323,1325,1327,1329,1331,1333,1335,1337,1339,1341,1343,1345,1347,1349,1351,1353,1355,1357,1359,1361,1363,1365,1367,1369,1371,1373,1375,1377,1379,1381,1383,1385,1387,1389,1391,1393,1395,1397,1399,1401,1403,1405,1407,1409,1411,1413,1415,1417,1419,1421,1423,1425,1427,1429,1431,1433,1435,1437,1439,1441,1443,1445,1447,1449,1451,1453,1455,1457,1459,1461,1463,1465,1467,1469,1471,1473,1475,1477,1479,1481,1483,1485,1487,1489,1491,1493,1495,1497,1499,1501,1503,1505,1507,1509,1511,1513,1515,1517,1519,1521,1523,1525,1527,1529,1531,1533,1535,1537,1539,1541,1543,1545,1547,1549,1551,1553,1555,1557,1559,1561,1563,1565,1567,1569,1571,1573,1575,1577,1579,1581,1583,1585,1587,1589,1591,1593,1595,1597,1599,1601,1603,1605,1607,1609,1611,1613,1615,1617,1619,1621,1623,1625,1627,1629,1631,1633,1635,1637,1639,1641,1643,1645,1647,1649,1651,1653,1655,1657,1659,1661,1663,1665,1667,1669,1671,1673,1675,1677,1679,1681,1683,1685,1687,1689,1691,1693,1695,1697,1699,1701,1703,1705,1707,1709,1711,1713,1715,1717,1719,1721,1723,1725,1727,1729,1731,1733,1735,1737,1739,1741,1743,1745,1747,1749,1751,1753,1755,1757,1759,1761,1763,1765,1767,1769,1771,1773,1775,1777,1779,1781,1783,1785,1787,1789,1791,1793,1795,1797,1799,1801,1803,1805,1807,1809,1811,1813,1815,1817,1819,1821,1823,1825,1827,1829,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,1831,1833,1835,1837,1839,1841,1843,1845,1847,1849,1851,1853,1855,1857,1859,1861,1863,1865,1867,1869,1871,1873,1875,1877,1879,1881,1883,1885,1887,1889,1891,1893,1895,1897,1899,1901,1903,1905,1907,1909,1911,1913,1915,1917,1919,1921,1923,1925,1927,1929,1931,1933,1935,1937,1939,1941,1943,1945,1947,1949,1951,1953,1955,1957,1959,1961,1963,1965,1967,1969,1971,1973,1975,1977,1979,1981,1983,1985,1987,1989,1991,1993,1995,1997,1999,2001,2003,2005,2007,2009,2011,2013,2015,2017,2019,2021,2023,2025,2027,2029,2031,2033,2035,2037,2039,2041,2043,2045,2047,2049,2051,2053,2055,2057,2059,2061,2063,2065,2067,2069,2071,2073,2075,2077,2079,2081,2083,2085,2087,2089,2091,2093,2095,2097,2099,2101,2103,2105,2107,2109,2111,2113,2115,2117,2119,2121,2123,2125,2127,2129,2131,2133,2135,2137,2139,2141,2143,2145,2147,2149,2151,2153,2155,2157,2159,2161,2163,2165,2167,2169,2171,2173,2175,2177,2179,2181,2183,2185,2187,2189,2191,2193,2195,2197,2199,2201,2203,2205,2207,2209,2211,2213,2215,2217,2219,2221,2223,2225,2227,2229,2231,2233,2235,2237,2239,2241,2243,2245,2247,2249,2251,2253,2255,2257,2259,2261,2263,2265,2267,2269,2271,2273,2275,2277,2279,2281,2283,2285,2287,2289,2291,2293,2295,2297,2299,2301,2303,2305,2307,2309,2311,2313,2315,2317,2319,2321,2323,2325,2327,2329,2331,2333,2335,2337,2339,2341,2343,2345,2347,2349,2351,2353,2355,2357,2359,2361,2363,2365,2367,2369,2371,2373,2375,2377,2379,2381,2383,2385,2387,2389,2391,2393,2395,2397,2399,2401,2403,2405,2407,2409,2411,2413,2415,2417,2419,2421,2423,2425,2427,2429,2431,2433,2435,2437,2439,2441,2443,2445,2447,2449,2451,2453,2455,2457,2459,2461,2463,2465,2467,2469,2471,2473,2475,2477,2479,2481,2483,2485,2487,2489,2491,2493,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,2495,2497,2499,2501,2503,2505,2507,2509,2511,2513,2515,2517,2519,2521,2523,2525,2527,2529,2531,2533,2535,2537,2539,2541,2543,2545,2547,2549,2551,2553,2555,2557,2559,2561,2563,2565,2567,2569,2571,2573,2575,2577,2579,2581,2583,2585,2587,2589,2591,2593,2595,2597,2599,2601,2603,2605,2607,2609,2611,2613,2615,2617,2619,2621,2623,2625,2627,2629,2631,2633,2635,2637,2639,2641,2643,2645,2647,2649,2651,2653,2655,2657,2659,2661,2663,2665,2667,2669,2671,2673,2675,2677,2679,2681,2683,2685,2687,2689,2691,2693,2695,2697,2699,2701,2703,2705,2707,2709,2711,2713,2715,2717,2719,2721,2723,2725,2727,2729,2731,2733,2735,2737,2739,2741,2743,2745,2747,2749,2751,2753,2755,2757,2759,2761,2763,2765,2767,2769,2771,2773,2775,2777,2779,2781,2783,2785,2787,2789,2791,2793,2795,2797,2799,2801,2803,2805,2807,2809,2811,2813,2815,2817,2819,2821,2823,2825,2827,2829,2831,2833,2835,2837,2839,2841,2843,2845,2847,2849,2851,2853,2855,2857,2859,2861,2863,2865,2867,2869,2871,2873,2875,2877,2879,2881,2883,2885,2887,2889,2891,2893,2895,2897,2899,2901,2903,2905,2907,2909,2911,2913,2915,2917,2919,2921,2923,2925,2927,2929,2931,2933,2935,2937,2939,2941,2943,2945,2947,2949,2951,2953,2955,2957,2959,2961,2963,2965,2967,2969,2971,2973,2975,2977,2979,2981,2983,2985,2987,2989,2991,2993,2995,2997,2999,3001,3003,3005,3007,3009,3011,3013,3015,3017,3019,3021,3023,3025,3027,3029,3031,3033,3035,3037,3039,3041,3043,3045,3047,3049,3051,3053,3055,3057,3059,3061,3063,3065,3067,3069,3071,3073,3075,3077,3079,3081,3083,3085,3087,3089,3091,3093,3095,3097,3099,3101,3103,3105,3107,3109,3111,3113,3115,3117,3119,3121,3123,3125,3127,3129,3131,3133,3135,3137,3139,3141,3143,3145,3147,3149,3151,3153,3155,3157,3159,3161,3163,3165,3167,3169,3171,3173,3175,3177,3179,3181,3183,3185,3187,3189,3191,3193,3195,3197,3199,3201,3203,3205,3207,3209,3211,3213,3215,3217,3219,3221,3223,3225,3227,3229,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,3231,3233,3235,3237,3239,3241,3243,3245,3247,3249,3251,3253,3255,3257,3259,3261,3263,3265,3267,3269,3271,3273,3275,3277,3279,3281,3283,3285,3287,3289,3291,3293,3295,3297,3299,3301,3303,3305,3307,3309,3311,3313,3315,3317,3319,3321,3323,3325,3327,3329,3331,3333,3335,3337,3339,3341,3343,3345,3347,3349,3351,3353,3355,3357,3359,3361,3363,3365,3367,3369,3371,3373,3375,3377,3379,3381,3383,3385,3387,3389,3391,3393,3395,3397,3399,3401,3403,3405,3407,3409,3411,3413,3415,3417,3419,3421,3423,3425,3427,3429,3431,3433,3435,3437,3439,3441,3443,3445,3447,3449,3451,3453,3455,3457,3459,3461,3463,3465,3467,3469,3471,3473,3475,3477,3479,3481,3483,3485,3487,3489,3491,3493,3495,3497,3499,3501,3503,3505,3507,3509,3511,3513,3515,3517,3519,3521,3523,3525,3527,3529,3531,3533,3535,3537,3539,3541,3543,3545,3547,3549,3551,3553,3555,3557,3559,3561,3563,3565,3567,3569,3571,3573,3575,3577,3579,3581,3583,3585,3587,3589,3591,3593,3595,3597,3599,3601,3603,3605,3607,3609,3611,3613,3615,3617,3619,3621,3623,3625,3627,3629,3631,3633,3635,3637,3639,3641,3643,3645,3647,3649,3651,3653,3655,3657,3659,3661,3663,3665,3667,3669,3671,3673,3675,3677,3679,3681,3683,3685,3687,3689,3691,3693,3695,3697,3699,3701,3703,3705,3707,3709,3711,3713,3715,3717,3719,3721,3723,3725,3727,3729,3731,3733,3735,3737,3739,3741,3743,3745,3747,3749,3751,3753,3755,3757,3759,3761,3763,3765,3767,3769,3771,3773,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,3775,3777,3779,3781,3783,3785,3787,3789,3791,3793,3795,3797,3799,3801,3803,3805,3807,3809,3811,3813,3815,3817,3819,3821,3823,3825,3827,3829,3831,3833,3835,3837,3839,3841,3843,3845,3847,3849,3851,3853,3855,3857,3859,3861,3863,3865,3867,3869,3871,3873,3875,3877,3879,3881,3883,3885,3887,3889,3891,3893,3895,3897,3899,3901,3903,3905,3907,3909,3911,3913,3915,3917,3919,3921,3923,3925,3927,3929,3931,3933,3935,3937,3939,3941,3943,3945,3947,3949,3951,3953,3955,3957,3959,3961,3963,3965,3967,3969,3971,3973,3975,3977,3979,3981,3983,3985,3987,3989,3991,3993,3995,3997,3999,4001,4003,4005,4007,4009,4011,4013,4015,4017,4019,4021,4023,4025,4027,4029,4031,4033,4035,4037,4039,4041,4043,4045,4047,4049,4051,4053,4055,4057,4059,4061,4063,4065,4067,4069,4071,4073,4075,4077,4079,4081,4083,4085,4087,4089,4091,4093,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1);
 constant children_right : intArray(nNodes-1 downto 0)  :=  (2,4,6,8,12,10,14,16,28,18,30,26,22,20,24,32,60,34,62,58,54,36,56,52,50,48,46,44,40,38,42,64,114,734,66,116,112,108,68,110,106,104,102,100,98,94,70,96,92,736,90,738,88,86,84,82,80,78,76,740,742,74,72,118,744,198,746,748,750,120,200,196,192,122,752,194,190,188,186,184,182,178,754,124,180,176,756,758,174,172,170,168,166,164,162,160,760,158,156,154,152,148,126,150,146,144,142,140,138,136,134,132,130,762,764,766,128,768,770,202,308,204,310,306,772,774,302,776,778,206,304,300,780,298,782,296,294,784,786,788,790,292,288,208,290,286,284,282,792,280,278,276,274,272,270,268,266,264,794,262,796,798,800,258,210,260,256,254,252,250,248,802,804,806,808,246,244,810,242,240,238,812,236,234,232,230,814,816,818,228,226,224,222,820,220,218,216,822,824,214,212,312,454,314,456,452,826,828,448,316,830,450,832,446,444,834,442,440,438,434,836,318,436,432,430,428,426,838,424,840,842,422,420,844,846,848,418,416,414,412,410,850,852,854,408,856,858,404,320,860,862,406,402,400,398,396,394,864,866,868,392,390,388,386,384,870,872,874,382,380,378,376,374,372,370,368,366,364,362,876,360,358,356,354,352,350,348,346,342,878,880,882,884,322,886,344,340,888,890,892,338,336,334,332,330,328,894,896,898,326,324,458,900,902,588,904,906,460,908,590,586,582,462,910,912,584,914,916,918,580,920,578,576,574,572,922,924,926,928,930,932,934,936,568,938,940,942,464,570,566,944,564,562,560,558,556,946,948,950,554,552,550,548,546,952,954,544,542,538,956,958,960,962,466,964,540,966,968,970,972,974,536,534,532,976,978,980,982,984,530,986,988,990,992,528,526,524,522,520,994,518,516,996,998,1000,514,1002,1004,1006,1008,1010,1012,1014,512,510,508,506,504,1016,502,500,498,496,1018,1020,494,492,1022,490,1024,488,1026,1028,486,1030,484,482,480,1032,476,1034,468,1036,478,474,472,1038,1040,1042,470,1044,1046,1048,1050,1052,1054,1056,592,1058,1060,730,1062,594,1064,732,1066,728,1068,1070,1072,1074,724,1076,596,726,722,1078,720,718,716,1080,1082,1084,714,710,1086,1088,1090,1092,1094,1096,598,712,1098,708,1100,1102,706,704,1104,702,1106,1108,1110,700,1112,1114,1116,698,696,1118,694,692,690,688,686,1120,684,680,600,682,678,676,674,1122,672,1124,670,1126,1128,668,666,1130,1132,664,1134,1136,1138,662,660,658,656,654,1140,1142,652,650,648,646,1144,644,1146,642,1148,1150,1152,640,638,636,1154,1156,634,632,630,628,626,624,1158,622,618,602,620,1160,1162,1164,1166,616,614,1168,612,1170,1172,1174,1176,1178,610,608,606,604,1180,1182,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,1184,1186,1188,1190,1192,1194,1196,1198,1200,1202,1204,1206,1208,1210,1212,1214,1216,1218,1220,1222,1224,1226,1228,1230,1232,1234,1236,1238,1240,1242,1244,1246,1248,1250,1252,1254,1256,1258,1260,1262,1264,1266,1268,1270,1272,1274,1276,1278,1280,1282,1284,1286,1288,1290,1292,1294,1296,1298,1300,1302,1304,1306,1308,1310,1312,1314,1316,1318,1320,1322,1324,1326,1328,1330,1332,1334,1336,1338,1340,1342,1344,1346,1348,1350,1352,1354,1356,1358,1360,1362,1364,1366,1368,1370,1372,1374,1376,1378,1380,1382,1384,1386,1388,1390,1392,1394,1396,1398,1400,1402,1404,1406,1408,1410,1412,1414,1416,1418,1420,1422,1424,1426,1428,1430,1432,1434,1436,1438,1440,1442,1444,1446,1448,1450,1452,1454,1456,1458,1460,1462,1464,1466,1468,1470,1472,1474,1476,1478,1480,1482,1484,1486,1488,1490,1492,1494,1496,1498,1500,1502,1504,1506,1508,1510,1512,1514,1516,1518,1520,1522,1524,1526,1528,1530,1532,1534,1536,1538,1540,1542,1544,1546,1548,1550,1552,1554,1556,1558,1560,1562,1564,1566,1568,1570,1572,1574,1576,1578,1580,1582,1584,1586,1588,1590,1592,1594,1596,1598,1600,1602,1604,1606,1608,1610,1612,1614,1616,1618,1620,1622,1624,1626,1628,1630,1632,1634,1636,1638,1640,1642,1644,1646,1648,1650,1652,1654,1656,1658,1660,1662,1664,1666,1668,1670,1672,1674,1676,1678,1680,1682,1684,1686,1688,1690,1692,1694,1696,1698,1700,1702,1704,1706,1708,1710,1712,1714,1716,1718,1720,1722,1724,1726,1728,1730,1732,1734,1736,1738,1740,1742,1744,1746,1748,1750,1752,1754,1756,1758,1760,1762,1764,1766,1768,1770,1772,1774,1776,1778,1780,1782,1784,1786,1788,1790,1792,1794,1796,1798,1800,1802,1804,1806,1808,1810,1812,1814,1816,1818,1820,1822,1824,1826,1828,1830,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,1832,1834,1836,1838,1840,1842,1844,1846,1848,1850,1852,1854,1856,1858,1860,1862,1864,1866,1868,1870,1872,1874,1876,1878,1880,1882,1884,1886,1888,1890,1892,1894,1896,1898,1900,1902,1904,1906,1908,1910,1912,1914,1916,1918,1920,1922,1924,1926,1928,1930,1932,1934,1936,1938,1940,1942,1944,1946,1948,1950,1952,1954,1956,1958,1960,1962,1964,1966,1968,1970,1972,1974,1976,1978,1980,1982,1984,1986,1988,1990,1992,1994,1996,1998,2000,2002,2004,2006,2008,2010,2012,2014,2016,2018,2020,2022,2024,2026,2028,2030,2032,2034,2036,2038,2040,2042,2044,2046,2048,2050,2052,2054,2056,2058,2060,2062,2064,2066,2068,2070,2072,2074,2076,2078,2080,2082,2084,2086,2088,2090,2092,2094,2096,2098,2100,2102,2104,2106,2108,2110,2112,2114,2116,2118,2120,2122,2124,2126,2128,2130,2132,2134,2136,2138,2140,2142,2144,2146,2148,2150,2152,2154,2156,2158,2160,2162,2164,2166,2168,2170,2172,2174,2176,2178,2180,2182,2184,2186,2188,2190,2192,2194,2196,2198,2200,2202,2204,2206,2208,2210,2212,2214,2216,2218,2220,2222,2224,2226,2228,2230,2232,2234,2236,2238,2240,2242,2244,2246,2248,2250,2252,2254,2256,2258,2260,2262,2264,2266,2268,2270,2272,2274,2276,2278,2280,2282,2284,2286,2288,2290,2292,2294,2296,2298,2300,2302,2304,2306,2308,2310,2312,2314,2316,2318,2320,2322,2324,2326,2328,2330,2332,2334,2336,2338,2340,2342,2344,2346,2348,2350,2352,2354,2356,2358,2360,2362,2364,2366,2368,2370,2372,2374,2376,2378,2380,2382,2384,2386,2388,2390,2392,2394,2396,2398,2400,2402,2404,2406,2408,2410,2412,2414,2416,2418,2420,2422,2424,2426,2428,2430,2432,2434,2436,2438,2440,2442,2444,2446,2448,2450,2452,2454,2456,2458,2460,2462,2464,2466,2468,2470,2472,2474,2476,2478,2480,2482,2484,2486,2488,2490,2492,2494,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,2496,2498,2500,2502,2504,2506,2508,2510,2512,2514,2516,2518,2520,2522,2524,2526,2528,2530,2532,2534,2536,2538,2540,2542,2544,2546,2548,2550,2552,2554,2556,2558,2560,2562,2564,2566,2568,2570,2572,2574,2576,2578,2580,2582,2584,2586,2588,2590,2592,2594,2596,2598,2600,2602,2604,2606,2608,2610,2612,2614,2616,2618,2620,2622,2624,2626,2628,2630,2632,2634,2636,2638,2640,2642,2644,2646,2648,2650,2652,2654,2656,2658,2660,2662,2664,2666,2668,2670,2672,2674,2676,2678,2680,2682,2684,2686,2688,2690,2692,2694,2696,2698,2700,2702,2704,2706,2708,2710,2712,2714,2716,2718,2720,2722,2724,2726,2728,2730,2732,2734,2736,2738,2740,2742,2744,2746,2748,2750,2752,2754,2756,2758,2760,2762,2764,2766,2768,2770,2772,2774,2776,2778,2780,2782,2784,2786,2788,2790,2792,2794,2796,2798,2800,2802,2804,2806,2808,2810,2812,2814,2816,2818,2820,2822,2824,2826,2828,2830,2832,2834,2836,2838,2840,2842,2844,2846,2848,2850,2852,2854,2856,2858,2860,2862,2864,2866,2868,2870,2872,2874,2876,2878,2880,2882,2884,2886,2888,2890,2892,2894,2896,2898,2900,2902,2904,2906,2908,2910,2912,2914,2916,2918,2920,2922,2924,2926,2928,2930,2932,2934,2936,2938,2940,2942,2944,2946,2948,2950,2952,2954,2956,2958,2960,2962,2964,2966,2968,2970,2972,2974,2976,2978,2980,2982,2984,2986,2988,2990,2992,2994,2996,2998,3000,3002,3004,3006,3008,3010,3012,3014,3016,3018,3020,3022,3024,3026,3028,3030,3032,3034,3036,3038,3040,3042,3044,3046,3048,3050,3052,3054,3056,3058,3060,3062,3064,3066,3068,3070,3072,3074,3076,3078,3080,3082,3084,3086,3088,3090,3092,3094,3096,3098,3100,3102,3104,3106,3108,3110,3112,3114,3116,3118,3120,3122,3124,3126,3128,3130,3132,3134,3136,3138,3140,3142,3144,3146,3148,3150,3152,3154,3156,3158,3160,3162,3164,3166,3168,3170,3172,3174,3176,3178,3180,3182,3184,3186,3188,3190,3192,3194,3196,3198,3200,3202,3204,3206,3208,3210,3212,3214,3216,3218,3220,3222,3224,3226,3228,3230,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,3232,3234,3236,3238,3240,3242,3244,3246,3248,3250,3252,3254,3256,3258,3260,3262,3264,3266,3268,3270,3272,3274,3276,3278,3280,3282,3284,3286,3288,3290,3292,3294,3296,3298,3300,3302,3304,3306,3308,3310,3312,3314,3316,3318,3320,3322,3324,3326,3328,3330,3332,3334,3336,3338,3340,3342,3344,3346,3348,3350,3352,3354,3356,3358,3360,3362,3364,3366,3368,3370,3372,3374,3376,3378,3380,3382,3384,3386,3388,3390,3392,3394,3396,3398,3400,3402,3404,3406,3408,3410,3412,3414,3416,3418,3420,3422,3424,3426,3428,3430,3432,3434,3436,3438,3440,3442,3444,3446,3448,3450,3452,3454,3456,3458,3460,3462,3464,3466,3468,3470,3472,3474,3476,3478,3480,3482,3484,3486,3488,3490,3492,3494,3496,3498,3500,3502,3504,3506,3508,3510,3512,3514,3516,3518,3520,3522,3524,3526,3528,3530,3532,3534,3536,3538,3540,3542,3544,3546,3548,3550,3552,3554,3556,3558,3560,3562,3564,3566,3568,3570,3572,3574,3576,3578,3580,3582,3584,3586,3588,3590,3592,3594,3596,3598,3600,3602,3604,3606,3608,3610,3612,3614,3616,3618,3620,3622,3624,3626,3628,3630,3632,3634,3636,3638,3640,3642,3644,3646,3648,3650,3652,3654,3656,3658,3660,3662,3664,3666,3668,3670,3672,3674,3676,3678,3680,3682,3684,3686,3688,3690,3692,3694,3696,3698,3700,3702,3704,3706,3708,3710,3712,3714,3716,3718,3720,3722,3724,3726,3728,3730,3732,3734,3736,3738,3740,3742,3744,3746,3748,3750,3752,3754,3756,3758,3760,3762,3764,3766,3768,3770,3772,3774,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,3776,3778,3780,3782,3784,3786,3788,3790,3792,3794,3796,3798,3800,3802,3804,3806,3808,3810,3812,3814,3816,3818,3820,3822,3824,3826,3828,3830,3832,3834,3836,3838,3840,3842,3844,3846,3848,3850,3852,3854,3856,3858,3860,3862,3864,3866,3868,3870,3872,3874,3876,3878,3880,3882,3884,3886,3888,3890,3892,3894,3896,3898,3900,3902,3904,3906,3908,3910,3912,3914,3916,3918,3920,3922,3924,3926,3928,3930,3932,3934,3936,3938,3940,3942,3944,3946,3948,3950,3952,3954,3956,3958,3960,3962,3964,3966,3968,3970,3972,3974,3976,3978,3980,3982,3984,3986,3988,3990,3992,3994,3996,3998,4000,4002,4004,4006,4008,4010,4012,4014,4016,4018,4020,4022,4024,4026,4028,4030,4032,4034,4036,4038,4040,4042,4044,4046,4048,4050,4052,4054,4056,4058,4060,4062,4064,4066,4068,4070,4072,4074,4076,4078,4080,4082,4084,4086,4088,4090,4092,4094,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1);
 constant value_int : intArray(nNodes-1 downto 0)  :=  (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,-15872,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,42496,0,-61952,0,0,0,0,0,0,0,-1187328,-90112,0,0,0,-18432,0,-22016,102912,-512,0,0,0,0,0,48128,0,0,0,0,0,0,0,-211968,0,0,0,103424,3072,0,0,0,0,0,0,0,0,22528,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,-65024,41472,51712,0,-667648,-64000,0,0,0,0,0,181760,-85504,0,-239616,-2048,0,0,0,-156160,0,-86528,0,0,-57344,62464,-416768,11264,0,0,0,0,0,0,0,8704,0,0,0,0,0,0,0,0,0,48128,0,-140800,-74752,11776,0,0,0,0,0,0,0,0,193536,-66560,195072,9728,0,0,-41984,0,0,0,-3584,0,0,0,0,-24576,23552,-102400,0,0,0,0,-37888,0,0,0,-28672,-583680,0,0,0,0,0,0,0,-172032,-43008,0,0,-30720,0,-15872,0,0,-33280,0,0,0,0,125952,0,0,0,0,0,0,-66560,0,93184,-3072,0,0,3072,-148992,33792,0,0,0,0,0,-22528,93184,75776,0,-241664,16896,0,0,-27648,110592,0,0,0,0,0,0,0,-86016,231936,0,0,0,0,0,48640,-133120,-74240,0,0,0,0,0,0,0,0,0,0,0,58880,0,0,0,0,0,0,0,0,0,-115200,26112,-28672,101376,0,6144,0,0,123904,-24576,-52224,0,0,0,0,0,0,-169984,75264,-69120,0,0,0,-11264,7168,0,-24064,-659456,0,-15872,0,0,0,0,25600,-76288,0,-13824,-31232,71680,0,6656,0,0,0,0,77312,-120832,115712,-17920,-107520,28672,10240,-325120,0,-512,-74752,88576,0,0,0,48640,0,0,0,0,0,16384,-37888,79360,0,0,0,0,0,32768,97792,0,0,0,13824,-44544,121856,-24064,0,-98304,0,-75264,-11776,90624,-127488,16896,0,0,0,4096,-20992,49664,30720,-54272,0,-26112,24064,-65024,-60416,0,0,0,0,0,32768,0,0,-68608,-9216,175616,0,67072,7680,-51200,-25088,246272,-2048,-83456,0,0,0,0,0,20992,0,0,0,0,-17920,76800,0,0,75264,0,29696,0,71168,-29696,0,-36352,0,0,0,31232,0,-97280,0,-9728,0,0,0,41984,288256,-14336,0,16384,-46592,106496,10240,-41984,-7168,18944,0,-9216,-4608,0,-17408,0,-142336,0,-40448,0,1024,165376,46080,691200,0,15360,0,0,0,-46592,0,0,0,-276992,-80896,9216,0,0,38400,-8192,-4096,-165888,-46592,26624,0,0,-5120,0,-11776,165888,0,0,-35840,0,31232,-72192,249344,0,14848,-95744,326656,0,0,108544,0,0,0,0,0,-36352,0,0,0,0,0,0,0,17408,0,66048,0,-15360,-143872,0,0,6656,-40960,0,-59904,-3584,42496,0,0,0,0,0,25600,-49664,0,0,0,0,14848,0,-119296,0,-16384,-320000,44032,0,0,0,-86016,37888,0,0,0,0,0,0,-33792,0,0,0,0,-25088,-68608,38912,86016,0,0,-40448,0,-8704,-71680,16896,-394752,-11776,0,0,0,0,224256,-15360,-823296,-77312,-550912,-137216,18944,258048,35840,455680,25600,-105472,-82432,112640,-141312,4608,-19968,20480,193536,1099776,16384,546816,68096,311808,-28160,158720,47616,-94208,-26624,203776,-21504,324096,-39936,-929792,-82432,59392,-201728,19968,-176128,8704,-99840,74240,7168,263680,58368,-82944,-30720,136704,2048,446464,71680,676352,109568,-41984,2048,-120320,-85504,48128,180736,8704,-23040,39424,-175104,-19968,31232,-270848,-49152,51712,-543744,-2560,-79872,59392,-82432,17920,229888,-17408,-202752,-2560,-23552,-726528,147456,2560,-43008,25088,19968,-174080,-300032,72704,-93696,124928,-500224,3072,118784,-41984,-78848,0,-19456,198144,-186880,29696,45568,-33280,67584,786944,-43008,76800,-53248,39936,-67072,80384,35328,742912,-12800,406016,-128512,23040,-21504,96256,3072,254976,-53760,25088,41472,-1536,137216,-26112,21504,-40448,-44032,-214528,-121344,24064,-18432,114176,-346112,4608,64000,-97280,64512,-9728,20992,273408,28672,-39424,-15872,-15872,42496,42496,-61952,-61952,-1187328,-1187328,-90112,-90112,-18432,-18432,-22016,-22016,102912,102912,-512,-512,48128,48128,-211968,-211968,103424,103424,3072,3072,22528,22528,-65024,-65024,41472,41472,51712,51712,-667648,-667648,-64000,-64000,181760,181760,-85504,-85504,-239616,-239616,-2048,-2048,-156160,-156160,-86528,-86528,-57344,-57344,62464,62464,-416768,-416768,11264,11264,8704,8704,48128,48128,-140800,-140800,-74752,-74752,11776,11776,193536,193536,-66560,-66560,195072,195072,9728,9728,-41984,-41984,-3584,-3584,-24576,-24576,23552,23552,-102400,-102400,-37888,-37888,-28672,-28672,-583680,-583680,-172032,-172032,-43008,-43008,-30720,-30720,-15872,-15872,-33280,-33280,125952,125952,-66560,-66560,93184,93184,-3072,-3072,3072,3072,-148992,-148992,33792,33792,-22528,-22528,93184,93184,75776,75776,-241664,-241664,16896,16896,-27648,-27648,110592,110592,0,0,-86016,-86016,231936,231936,48640,48640,-133120,-133120,-74240,-74240,58880,58880,-115200,-115200,26112,26112,-28672,-28672,101376,101376,6144,6144,123904,123904,-24576,-24576,-52224,-52224,-169984,-169984,75264,75264,-69120,-69120,-11264,-11264,7168,7168,-24064,-24064,-659456,-659456,-15872,-15872,25600,25600,-76288,-76288,-13824,-13824,-31232,-31232,71680,71680,6656,6656,77312,77312,-120832,-120832,115712,115712,-17920,-17920,-107520,-107520,28672,28672,10240,10240,-325120,-325120,-512,-512,-74752,-74752,88576,88576,48640,48640,16384,16384,-37888,-37888,79360,79360,32768,32768,97792,97792,13824,13824,-44544,-44544,121856,121856,-24064,-24064,-98304,-98304,-75264,-75264,-11776,-11776,90624,90624,-127488,-127488,16896,16896,4096,4096,-20992,-20992,49664,49664,30720,30720,-54272,-54272,-26112,-26112,24064,24064,-65024,-65024,-60416,-60416,32768,32768,-68608,-68608,-9216,-9216,175616,175616,67072,67072,7680,7680,-51200,-51200,-25088,-25088,246272,246272,-2048,-2048,-83456,-83456,20992,20992,-17920,-17920,76800,76800,75264,75264,29696,29696,71168,71168,-29696,-29696,-36352,-36352,31232,31232,-97280,-97280,-9728,-9728,41984,41984,288256,288256,-14336,-14336,16384,16384,-46592,-46592,106496,106496,10240,10240,-41984,-41984,-7168,-7168,18944,18944,-9216,-9216,-4608,-4608,-17408,-17408,-142336,-142336,-40448,-40448,1024,1024,165376,165376,46080,46080,691200,691200,15360,15360,-46592,-46592,-276992,-276992,-80896,-80896,9216,9216,38400,38400,-8192,-8192,-4096,-4096,-165888,-165888,-46592,-46592,26624,26624,-5120,-5120,-11776,-11776,165888,165888,-35840,-35840,31232,31232,-72192,-72192,249344,249344,14848,14848,-95744,-95744,326656,326656,108544,108544,-36352,-36352,17408,17408,66048,66048,-15360,-15360,-143872,-143872,6656,6656,-40960,-40960,-59904,-59904,-3584,-3584,42496,42496,25600,25600,-49664,-49664,14848,14848,-119296,-119296,-16384,-16384,-320000,-320000,44032,44032,-86016,-86016,37888,37888,-33792,-33792,-25088,-25088,-68608,-68608,38912,38912,86016,86016,-40448,-40448,-8704,-8704,-71680,-71680,16896,16896,-394752,-394752,-11776,-11776,224256,224256,-15360,-15360,-15872,-15872,-15872,-15872,42496,42496,42496,42496,-61952,-61952,-61952,-61952,-1187328,-1187328,-1187328,-1187328,-90112,-90112,-90112,-90112,-18432,-18432,-18432,-18432,-22016,-22016,-22016,-22016,102912,102912,102912,102912,-512,-512,-512,-512,48128,48128,48128,48128,-211968,-211968,-211968,-211968,103424,103424,103424,103424,3072,3072,3072,3072,22528,22528,22528,22528,-65024,-65024,-65024,-65024,41472,41472,41472,41472,51712,51712,51712,51712,-667648,-667648,-667648,-667648,-64000,-64000,-64000,-64000,181760,181760,181760,181760,-85504,-85504,-85504,-85504,-239616,-239616,-239616,-239616,-2048,-2048,-2048,-2048,-156160,-156160,-156160,-156160,-86528,-86528,-86528,-86528,-57344,-57344,-57344,-57344,62464,62464,62464,62464,-416768,-416768,-416768,-416768,11264,11264,11264,11264,8704,8704,8704,8704,48128,48128,48128,48128,-140800,-140800,-140800,-140800,-74752,-74752,-74752,-74752,11776,11776,11776,11776,193536,193536,193536,193536,-66560,-66560,-66560,-66560,195072,195072,195072,195072,9728,9728,9728,9728,-41984,-41984,-41984,-41984,-3584,-3584,-3584,-3584,-24576,-24576,-24576,-24576,23552,23552,23552,23552,-102400,-102400,-102400,-102400,-37888,-37888,-37888,-37888,-28672,-28672,-28672,-28672,-583680,-583680,-583680,-583680,-172032,-172032,-172032,-172032,-43008,-43008,-43008,-43008,-30720,-30720,-30720,-30720,-15872,-15872,-15872,-15872,-33280,-33280,-33280,-33280,125952,125952,125952,125952,-66560,-66560,-66560,-66560,93184,93184,93184,93184,-3072,-3072,-3072,-3072,3072,3072,3072,3072,-148992,-148992,-148992,-148992,33792,33792,33792,33792,-22528,-22528,-22528,-22528,93184,93184,93184,93184,75776,75776,75776,75776,-241664,-241664,-241664,-241664,16896,16896,16896,16896,-27648,-27648,-27648,-27648,110592,110592,110592,110592,0,0,0,0,-86016,-86016,-86016,-86016,231936,231936,231936,231936,48640,48640,48640,48640,-133120,-133120,-133120,-133120,-74240,-74240,-74240,-74240,58880,58880,58880,58880,-115200,-115200,-115200,-115200,26112,26112,26112,26112,-28672,-28672,-28672,-28672,101376,101376,101376,101376,6144,6144,6144,6144,123904,123904,123904,123904,-24576,-24576,-24576,-24576,-52224,-52224,-52224,-52224,-169984,-169984,-169984,-169984,75264,75264,75264,75264,-69120,-69120,-69120,-69120,-11264,-11264,-11264,-11264,7168,7168,7168,7168,-24064,-24064,-24064,-24064,-659456,-659456,-659456,-659456,-15872,-15872,-15872,-15872,25600,25600,25600,25600,-76288,-76288,-76288,-76288,-13824,-13824,-13824,-13824,-31232,-31232,-31232,-31232,71680,71680,71680,71680,6656,6656,6656,6656,77312,77312,77312,77312,-120832,-120832,-120832,-120832,115712,115712,115712,115712,-17920,-17920,-17920,-17920,-107520,-107520,-107520,-107520,28672,28672,28672,28672,10240,10240,10240,10240,-325120,-325120,-325120,-325120,-512,-512,-512,-512,-74752,-74752,-74752,-74752,88576,88576,88576,88576,48640,48640,48640,48640,16384,16384,16384,16384,-37888,-37888,-37888,-37888,79360,79360,79360,79360,32768,32768,32768,32768,97792,97792,97792,97792,13824,13824,13824,13824,-44544,-44544,-44544,-44544,121856,121856,121856,121856,-24064,-24064,-24064,-24064,-98304,-98304,-98304,-98304,-75264,-75264,-75264,-75264,-11776,-11776,-11776,-11776,90624,90624,90624,90624,-127488,-127488,-127488,-127488,16896,16896,16896,16896,4096,4096,4096,4096,-20992,-20992,-20992,-20992,49664,49664,49664,49664,30720,30720,30720,30720,-54272,-54272,-54272,-54272,-26112,-26112,-26112,-26112,24064,24064,24064,24064,-65024,-65024,-65024,-65024,-60416,-60416,-60416,-60416,32768,32768,32768,32768,-68608,-68608,-68608,-68608,-9216,-9216,-9216,-9216,175616,175616,175616,175616,67072,67072,67072,67072,7680,7680,7680,7680,-51200,-51200,-51200,-51200,-25088,-25088,-25088,-25088,246272,246272,246272,246272,-2048,-2048,-2048,-2048,-83456,-83456,-83456,-83456,20992,20992,20992,20992,-17920,-17920,-17920,-17920,76800,76800,76800,76800,75264,75264,75264,75264,29696,29696,29696,29696,71168,71168,71168,71168,-29696,-29696,-29696,-29696,-36352,-36352,-36352,-36352,31232,31232,31232,31232,-97280,-97280,-97280,-97280,-9728,-9728,-9728,-9728,41984,41984,41984,41984,288256,288256,288256,288256,-14336,-14336,-14336,-14336,16384,16384,16384,16384,-46592,-46592,-46592,-46592,106496,106496,106496,106496,10240,10240,10240,10240,-41984,-41984,-41984,-41984,-7168,-7168,-7168,-7168,18944,18944,18944,18944,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,42496,42496,42496,42496,42496,42496,42496,42496,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,102912,102912,102912,102912,102912,102912,102912,102912,-512,-512,-512,-512,-512,-512,-512,-512,48128,48128,48128,48128,48128,48128,48128,48128,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,103424,103424,103424,103424,103424,103424,103424,103424,3072,3072,3072,3072,3072,3072,3072,3072,22528,22528,22528,22528,22528,22528,22528,22528,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,41472,41472,41472,41472,41472,41472,41472,41472,51712,51712,51712,51712,51712,51712,51712,51712,-667648,-667648,-667648,-667648,-667648,-667648,-667648,-667648,-64000,-64000,-64000,-64000,-64000,-64000,-64000,-64000,181760,181760,181760,181760,181760,181760,181760,181760,-85504,-85504,-85504,-85504,-85504,-85504,-85504,-85504,-239616,-239616,-239616,-239616,-239616,-239616,-239616,-239616,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-156160,-156160,-156160,-156160,-156160,-156160,-156160,-156160,-86528,-86528,-86528,-86528,-86528,-86528,-86528,-86528,-57344,-57344,-57344,-57344,-57344,-57344,-57344,-57344,62464,62464,62464,62464,62464,62464,62464,62464,-416768,-416768,-416768,-416768,-416768,-416768,-416768,-416768,11264,11264,11264,11264,11264,11264,11264,11264,8704,8704,8704,8704,8704,8704,8704,8704,48128,48128,48128,48128,48128,48128,48128,48128,-140800,-140800,-140800,-140800,-140800,-140800,-140800,-140800,-74752,-74752,-74752,-74752,-74752,-74752,-74752,-74752,11776,11776,11776,11776,11776,11776,11776,11776,193536,193536,193536,193536,193536,193536,193536,193536,-66560,-66560,-66560,-66560,-66560,-66560,-66560,-66560,195072,195072,195072,195072,195072,195072,195072,195072,9728,9728,9728,9728,9728,9728,9728,9728,-41984,-41984,-41984,-41984,-41984,-41984,-41984,-41984,-3584,-3584,-3584,-3584,-3584,-3584,-3584,-3584,-24576,-24576,-24576,-24576,-24576,-24576,-24576,-24576,23552,23552,23552,23552,23552,23552,23552,23552,-102400,-102400,-102400,-102400,-102400,-102400,-102400,-102400,-37888,-37888,-37888,-37888,-37888,-37888,-37888,-37888,-28672,-28672,-28672,-28672,-28672,-28672,-28672,-28672,-583680,-583680,-583680,-583680,-583680,-583680,-583680,-583680,-172032,-172032,-172032,-172032,-172032,-172032,-172032,-172032,-43008,-43008,-43008,-43008,-43008,-43008,-43008,-43008,-30720,-30720,-30720,-30720,-30720,-30720,-30720,-30720,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-33280,-33280,-33280,-33280,-33280,-33280,-33280,-33280,125952,125952,125952,125952,125952,125952,125952,125952,-66560,-66560,-66560,-66560,-66560,-66560,-66560,-66560,93184,93184,93184,93184,93184,93184,93184,93184,-3072,-3072,-3072,-3072,-3072,-3072,-3072,-3072,3072,3072,3072,3072,3072,3072,3072,3072,-148992,-148992,-148992,-148992,-148992,-148992,-148992,-148992,33792,33792,33792,33792,33792,33792,33792,33792,-22528,-22528,-22528,-22528,-22528,-22528,-22528,-22528,93184,93184,93184,93184,93184,93184,93184,93184,75776,75776,75776,75776,75776,75776,75776,75776,-241664,-241664,-241664,-241664,-241664,-241664,-241664,-241664,16896,16896,16896,16896,16896,16896,16896,16896,-27648,-27648,-27648,-27648,-27648,-27648,-27648,-27648,110592,110592,110592,110592,110592,110592,110592,110592,0,0,0,0,0,0,0,0,-86016,-86016,-86016,-86016,-86016,-86016,-86016,-86016,231936,231936,231936,231936,231936,231936,231936,231936,48640,48640,48640,48640,48640,48640,48640,48640,-133120,-133120,-133120,-133120,-133120,-133120,-133120,-133120,-74240,-74240,-74240,-74240,-74240,-74240,-74240,-74240,58880,58880,58880,58880,58880,58880,58880,58880,-115200,-115200,-115200,-115200,-115200,-115200,-115200,-115200,26112,26112,26112,26112,26112,26112,26112,26112,-28672,-28672,-28672,-28672,-28672,-28672,-28672,-28672,101376,101376,101376,101376,101376,101376,101376,101376,6144,6144,6144,6144,6144,6144,6144,6144,123904,123904,123904,123904,123904,123904,123904,123904,-24576,-24576,-24576,-24576,-24576,-24576,-24576,-24576,-52224,-52224,-52224,-52224,-52224,-52224,-52224,-52224,-169984,-169984,-169984,-169984,-169984,-169984,-169984,-169984,75264,75264,75264,75264,75264,75264,75264,75264,-69120,-69120,-69120,-69120,-69120,-69120,-69120,-69120,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,102912,102912,102912,102912,102912,102912,102912,102912,102912,102912,102912,102912,102912,102912,102912,102912,-512,-512,-512,-512,-512,-512,-512,-512,-512,-512,-512,-512,-512,-512,-512,-512,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,103424,103424,103424,103424,103424,103424,103424,103424,103424,103424,103424,103424,103424,103424,103424,103424,3072,3072,3072,3072,3072,3072,3072,3072,3072,3072,3072,3072,3072,3072,3072,3072,22528,22528,22528,22528,22528,22528,22528,22528,22528,22528,22528,22528,22528,22528,22528,22528,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,41472,41472,41472,41472,41472,41472,41472,41472,41472,41472,41472,41472,41472,41472,41472,41472,51712,51712,51712,51712,51712,51712,51712,51712,51712,51712,51712,51712,51712,51712,51712,51712,-667648,-667648,-667648,-667648,-667648,-667648,-667648,-667648,-667648,-667648,-667648,-667648,-667648,-667648,-667648,-667648,-64000,-64000,-64000,-64000,-64000,-64000,-64000,-64000,-64000,-64000,-64000,-64000,-64000,-64000,-64000,-64000,181760,181760,181760,181760,181760,181760,181760,181760,181760,181760,181760,181760,181760,181760,181760,181760,-85504,-85504,-85504,-85504,-85504,-85504,-85504,-85504,-85504,-85504,-85504,-85504,-85504,-85504,-85504,-85504,-239616,-239616,-239616,-239616,-239616,-239616,-239616,-239616,-239616,-239616,-239616,-239616,-239616,-239616,-239616,-239616,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-2048,-156160,-156160,-156160,-156160,-156160,-156160,-156160,-156160,-156160,-156160,-156160,-156160,-156160,-156160,-156160,-156160,-86528,-86528,-86528,-86528,-86528,-86528,-86528,-86528,-86528,-86528,-86528,-86528,-86528,-86528,-86528,-86528,-57344,-57344,-57344,-57344,-57344,-57344,-57344,-57344,-57344,-57344,-57344,-57344,-57344,-57344,-57344,-57344,62464,62464,62464,62464,62464,62464,62464,62464,62464,62464,62464,62464,62464,62464,62464,62464,-416768,-416768,-416768,-416768,-416768,-416768,-416768,-416768,-416768,-416768,-416768,-416768,-416768,-416768,-416768,-416768,11264,11264,11264,11264,11264,11264,11264,11264,11264,11264,11264,11264,11264,11264,11264,11264,8704,8704,8704,8704,8704,8704,8704,8704,8704,8704,8704,8704,8704,8704,8704,8704,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,-140800,-140800,-140800,-140800,-140800,-140800,-140800,-140800,-140800,-140800,-140800,-140800,-140800,-140800,-140800,-140800,-74752,-74752,-74752,-74752,-74752,-74752,-74752,-74752,-74752,-74752,-74752,-74752,-74752,-74752,-74752,-74752,11776,11776,11776,11776,11776,11776,11776,11776,11776,11776,11776,11776,11776,11776,11776,11776,193536,193536,193536,193536,193536,193536,193536,193536,193536,193536,193536,193536,193536,193536,193536,193536,-66560,-66560,-66560,-66560,-66560,-66560,-66560,-66560,-66560,-66560,-66560,-66560,-66560,-66560,-66560,-66560,195072,195072,195072,195072,195072,195072,195072,195072,195072,195072,195072,195072,195072,195072,195072,195072,9728,9728,9728,9728,9728,9728,9728,9728,9728,9728,9728,9728,9728,9728,9728,9728,-41984,-41984,-41984,-41984,-41984,-41984,-41984,-41984,-41984,-41984,-41984,-41984,-41984,-41984,-41984,-41984,-3584,-3584,-3584,-3584,-3584,-3584,-3584,-3584,-3584,-3584,-3584,-3584,-3584,-3584,-3584,-3584,-24576,-24576,-24576,-24576,-24576,-24576,-24576,-24576,-24576,-24576,-24576,-24576,-24576,-24576,-24576,-24576,23552,23552,23552,23552,23552,23552,23552,23552,23552,23552,23552,23552,23552,23552,23552,23552,-102400,-102400,-102400,-102400,-102400,-102400,-102400,-102400,-102400,-102400,-102400,-102400,-102400,-102400,-102400,-102400,-37888,-37888,-37888,-37888,-37888,-37888,-37888,-37888,-37888,-37888,-37888,-37888,-37888,-37888,-37888,-37888,-28672,-28672,-28672,-28672,-28672,-28672,-28672,-28672,-28672,-28672,-28672,-28672,-28672,-28672,-28672,-28672,-583680,-583680,-583680,-583680,-583680,-583680,-583680,-583680,-583680,-583680,-583680,-583680,-583680,-583680,-583680,-583680,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-18432,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,-22016,102912,102912,102912,102912,102912,102912,102912,102912,102912,102912,102912,102912,102912,102912,102912,102912,102912,102912,102912,102912,102912,102912,102912,102912,102912,102912,102912,102912,102912,102912,102912,102912,-512,-512,-512,-512,-512,-512,-512,-512,-512,-512,-512,-512,-512,-512,-512,-512,-512,-512,-512,-512,-512,-512,-512,-512,-512,-512,-512,-512,-512,-512,-512,-512,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,48128,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,-211968,103424,103424,103424,103424,103424,103424,103424,103424,103424,103424,103424,103424,103424,103424,103424,103424,103424,103424,103424,103424,103424,103424,103424,103424,103424,103424,103424,103424,103424,103424,103424,103424,3072,3072,3072,3072,3072,3072,3072,3072,3072,3072,3072,3072,3072,3072,3072,3072,3072,3072,3072,3072,3072,3072,3072,3072,3072,3072,3072,3072,3072,3072,3072,3072,22528,22528,22528,22528,22528,22528,22528,22528,22528,22528,22528,22528,22528,22528,22528,22528,22528,22528,22528,22528,22528,22528,22528,22528,22528,22528,22528,22528,22528,22528,22528,22528,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,-65024,41472,41472,41472,41472,41472,41472,41472,41472,41472,41472,41472,41472,41472,41472,41472,41472,41472,41472,41472,41472,41472,41472,41472,41472,41472,41472,41472,41472,41472,41472,41472,41472,51712,51712,51712,51712,51712,51712,51712,51712,51712,51712,51712,51712,51712,51712,51712,51712,51712,51712,51712,51712,51712,51712,51712,51712,51712,51712,51712,51712,51712,51712,51712,51712,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,-15872,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,42496,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-61952,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-1187328,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112,-90112);
 constant parent : intArray(nNodes-1 downto 0)  :=  (-1,0,0,1,1,2,2,3,3,5,5,4,4,6,6,7,7,9,9,13,13,12,12,14,14,11,11,8,8,10,10,15,15,17,17,21,21,29,29,28,28,30,30,27,27,26,26,25,25,24,24,23,23,20,20,22,22,19,19,16,16,18,18,31,31,34,34,38,38,46,46,62,62,61,61,58,58,57,57,56,56,55,55,54,54,53,53,52,52,50,50,48,48,45,45,47,47,44,44,43,43,42,42,41,41,40,40,37,37,39,39,36,36,32,32,35,35,63,63,69,69,73,73,83,83,102,102,116,116,112,112,111,111,110,110,109,109,108,108,107,107,106,106,105,105,104,104,101,101,103,103,100,100,99,99,98,98,97,97,95,95,94,94,93,93,92,92,91,91,90,90,89,89,88,88,85,85,81,81,84,84,80,80,79,79,78,78,77,77,76,76,72,72,75,75,71,71,65,65,70,70,119,119,121,121,129,129,143,143,164,164,200,200,199,199,196,196,195,195,194,194,192,192,191,191,190,190,189,189,185,185,184,184,183,183,182,182,180,180,179,179,178,178,176,176,175,175,170,170,169,169,168,168,167,167,166,166,163,163,165,165,159,159,157,157,156,156,155,155,154,154,153,153,152,152,151,151,150,150,149,149,147,147,146,146,145,145,142,142,144,144,141,141,136,136,135,135,133,133,131,131,126,126,130,130,123,123,120,120,122,122,201,201,203,203,209,209,221,221,248,248,293,293,310,310,309,309,305,305,304,304,303,303,302,302,301,301,300,300,296,296,288,288,295,295,287,287,286,286,285,285,284,284,283,283,282,282,281,281,280,280,278,278,277,277,276,276,275,275,274,274,273,273,272,272,271,271,270,270,269,269,268,268,264,264,263,263,262,262,261,261,260,260,256,256,255,255,254,254,253,253,252,252,247,247,251,251,244,244,240,240,239,239,238,238,237,237,236,236,232,232,231,231,228,228,226,226,225,225,224,224,223,223,219,219,222,222,218,218,217,217,216,216,214,214,213,213,208,208,211,211,205,205,202,202,204,204,311,311,317,317,322,322,347,347,373,373,441,441,449,449,445,445,444,444,439,439,443,443,437,437,436,436,435,435,433,433,430,430,428,428,426,426,425,425,422,422,421,421,420,420,419,419,417,417,416,416,415,415,414,414,413,413,405,405,401,401,400,400,398,398,397,397,396,396,395,395,394,394,389,389,383,383,382,382,381,381,368,368,375,375,367,367,366,366,363,363,362,362,361,361,360,360,359,359,355,355,354,354,353,353,352,352,351,351,349,349,343,343,348,348,334,334,333,333,332,332,331,331,329,329,321,321,325,325,320,320,314,314,319,319,457,457,462,462,473,473,491,491,519,519,570,570,588,588,587,587,586,586,585,585,579,579,577,577,576,576,569,569,571,571,568,568,566,566,565,565,564,564,563,563,562,562,561,561,558,558,557,557,556,556,552,552,550,550,548,548,547,547,546,546,545,545,542,542,541,541,540,540,539,539,538,538,534,534,531,531,530,530,527,527,525,525,523,523,522,522,521,521,518,518,520,520,517,517,515,515,514,514,513,513,512,512,511,511,509,509,508,508,504,504,500,500,498,498,497,497,494,494,484,484,492,492,483,483,479,479,478,478,477,477,475,475,471,471,474,474,466,466,460,460,464,464,33,33,49,49,51,51,59,59,60,60,64,64,66,66,67,67,68,68,74,74,82,82,86,86,87,87,96,96,113,113,114,114,115,115,117,117,118,118,124,124,125,125,127,127,128,128,132,132,134,134,137,137,138,138,139,139,140,140,148,148,158,158,160,160,161,161,162,162,171,171,172,172,173,173,174,174,177,177,181,181,186,186,187,187,188,188,193,193,197,197,198,198,206,206,207,207,210,210,212,212,215,215,220,220,227,227,229,229,230,230,233,233,234,234,235,235,241,241,242,242,243,243,245,245,246,246,249,249,250,250,257,257,258,258,259,259,265,265,266,266,267,267,279,279,289,289,290,290,291,291,292,292,294,294,297,297,298,298,299,299,306,306,307,307,308,308,312,312,313,313,315,315,316,316,318,318,323,323,324,324,326,326,327,327,328,328,330,330,335,335,336,336,337,337,338,338,339,339,340,340,341,341,342,342,344,344,345,345,346,346,350,350,356,356,357,357,358,358,364,364,365,365,369,369,370,370,371,371,372,372,374,374,376,376,377,377,378,378,379,379,380,380,384,384,385,385,386,386,387,387,388,388,390,390,391,391,392,392,393,393,399,399,402,402,403,403,404,404,406,406,407,407,408,408,409,409,410,410,411,411,412,412,418,418,423,423,424,424,427,427,429,429,431,431,432,432,434,434,438,438,440,440,442,442,446,446,447,447,448,448,450,450,451,451,452,452,453,453,454,454,455,455,456,456,458,458,459,459,461,461,463,463,465,465,467,467,468,468,469,469,470,470,472,472,476,476,480,480,481,481,482,482,485,485,486,486,487,487,488,488,489,489,490,490,493,493,495,495,496,496,499,499,501,501,502,502,503,503,505,505,506,506,507,507,510,510,516,516,524,524,526,526,528,528,529,529,532,532,533,533,535,535,536,536,537,537,543,543,544,544,549,549,551,551,553,553,554,554,555,555,559,559,560,560,567,567,572,572,573,573,574,574,575,575,578,578,580,580,581,581,582,582,583,583,584,584,589,589,590,590,733,733,734,734,735,735,736,736,737,737,738,738,739,739,740,740,741,741,742,742,743,743,744,744,745,745,746,746,747,747,748,748,749,749,750,750,751,751,752,752,753,753,754,754,755,755,756,756,757,757,758,758,759,759,760,760,761,761,762,762,763,763,764,764,765,765,766,766,767,767,768,768,769,769,770,770,771,771,772,772,773,773,774,774,775,775,776,776,777,777,778,778,779,779,780,780,781,781,782,782,783,783,784,784,785,785,786,786,787,787,788,788,789,789,790,790,791,791,792,792,793,793,794,794,795,795,796,796,797,797,798,798,799,799,800,800,801,801,802,802,803,803,804,804,805,805,806,806,807,807,808,808,809,809,810,810,811,811,812,812,813,813,814,814,815,815,816,816,817,817,818,818,819,819,820,820,821,821,822,822,823,823,824,824,825,825,826,826,827,827,828,828,829,829,830,830,831,831,832,832,833,833,834,834,835,835,836,836,837,837,838,838,839,839,840,840,841,841,842,842,843,843,844,844,845,845,846,846,847,847,848,848,849,849,850,850,851,851,852,852,853,853,854,854,855,855,856,856,857,857,858,858,859,859,860,860,861,861,862,862,863,863,864,864,865,865,866,866,867,867,868,868,869,869,870,870,871,871,872,872,873,873,874,874,875,875,876,876,877,877,878,878,879,879,880,880,881,881,882,882,883,883,884,884,885,885,886,886,887,887,888,888,889,889,890,890,891,891,892,892,893,893,894,894,895,895,896,896,897,897,898,898,899,899,900,900,901,901,902,902,903,903,904,904,905,905,906,906,907,907,908,908,909,909,910,910,911,911,912,912,913,913,914,914,915,915,916,916,917,917,918,918,919,919,920,920,921,921,922,922,923,923,924,924,925,925,926,926,927,927,928,928,929,929,930,930,931,931,932,932,933,933,934,934,935,935,936,936,937,937,938,938,939,939,940,940,941,941,942,942,943,943,944,944,945,945,946,946,947,947,948,948,949,949,950,950,951,951,952,952,953,953,954,954,955,955,956,956,957,957,958,958,959,959,960,960,961,961,962,962,963,963,964,964,965,965,966,966,967,967,968,968,969,969,970,970,971,971,972,972,973,973,974,974,975,975,976,976,977,977,978,978,979,979,980,980,981,981,982,982,983,983,984,984,985,985,986,986,987,987,988,988,989,989,990,990,991,991,992,992,993,993,994,994,995,995,996,996,997,997,998,998,999,999,1000,1000,1001,1001,1002,1002,1003,1003,1004,1004,1005,1005,1006,1006,1007,1007,1008,1008,1009,1009,1010,1010,1011,1011,1012,1012,1013,1013,1014,1014,1015,1015,1016,1016,1017,1017,1018,1018,1019,1019,1020,1020,1021,1021,1022,1022,1023,1023,1024,1024,1025,1025,1026,1026,1027,1027,1028,1028,1029,1029,1030,1030,1031,1031,1032,1032,1033,1033,1034,1034,1035,1035,1036,1036,1037,1037,1038,1038,1039,1039,1040,1040,1041,1041,1042,1042,1043,1043,1044,1044,1045,1045,1046,1046,1047,1047,1048,1048,1049,1049,1050,1050,1051,1051,1052,1052,1053,1053,1054,1054,1055,1055,1056,1056,1183,1183,1184,1184,1185,1185,1186,1186,1187,1187,1188,1188,1189,1189,1190,1190,1191,1191,1192,1192,1193,1193,1194,1194,1195,1195,1196,1196,1197,1197,1198,1198,1199,1199,1200,1200,1201,1201,1202,1202,1203,1203,1204,1204,1205,1205,1206,1206,1207,1207,1208,1208,1209,1209,1210,1210,1211,1211,1212,1212,1213,1213,1214,1214,1215,1215,1216,1216,1217,1217,1218,1218,1219,1219,1220,1220,1221,1221,1222,1222,1223,1223,1224,1224,1225,1225,1226,1226,1227,1227,1228,1228,1229,1229,1230,1230,1231,1231,1232,1232,1233,1233,1234,1234,1235,1235,1236,1236,1237,1237,1238,1238,1239,1239,1240,1240,1241,1241,1242,1242,1243,1243,1244,1244,1245,1245,1246,1246,1247,1247,1248,1248,1249,1249,1250,1250,1251,1251,1252,1252,1253,1253,1254,1254,1255,1255,1256,1256,1257,1257,1258,1258,1259,1259,1260,1260,1261,1261,1262,1262,1263,1263,1264,1264,1265,1265,1266,1266,1267,1267,1268,1268,1269,1269,1270,1270,1271,1271,1272,1272,1273,1273,1274,1274,1275,1275,1276,1276,1277,1277,1278,1278,1279,1279,1280,1280,1281,1281,1282,1282,1283,1283,1284,1284,1285,1285,1286,1286,1287,1287,1288,1288,1289,1289,1290,1290,1291,1291,1292,1292,1293,1293,1294,1294,1295,1295,1296,1296,1297,1297,1298,1298,1299,1299,1300,1300,1301,1301,1302,1302,1303,1303,1304,1304,1305,1305,1306,1306,1307,1307,1308,1308,1309,1309,1310,1310,1311,1311,1312,1312,1313,1313,1314,1314,1315,1315,1316,1316,1317,1317,1318,1318,1319,1319,1320,1320,1321,1321,1322,1322,1323,1323,1324,1324,1325,1325,1326,1326,1327,1327,1328,1328,1329,1329,1330,1330,1331,1331,1332,1332,1333,1333,1334,1334,1335,1335,1336,1336,1337,1337,1338,1338,1339,1339,1340,1340,1341,1341,1342,1342,1343,1343,1344,1344,1345,1345,1346,1346,1347,1347,1348,1348,1349,1349,1350,1350,1351,1351,1352,1352,1353,1353,1354,1354,1355,1355,1356,1356,1357,1357,1358,1358,1359,1359,1360,1360,1361,1361,1362,1362,1363,1363,1364,1364,1365,1365,1366,1366,1367,1367,1368,1368,1369,1369,1370,1370,1371,1371,1372,1372,1373,1373,1374,1374,1375,1375,1376,1376,1377,1377,1378,1378,1379,1379,1380,1380,1381,1381,1382,1382,1383,1383,1384,1384,1385,1385,1386,1386,1387,1387,1388,1388,1389,1389,1390,1390,1391,1391,1392,1392,1393,1393,1394,1394,1395,1395,1396,1396,1397,1397,1398,1398,1399,1399,1400,1400,1401,1401,1402,1402,1403,1403,1404,1404,1405,1405,1406,1406,1407,1407,1408,1408,1409,1409,1410,1410,1411,1411,1412,1412,1413,1413,1414,1414,1415,1415,1416,1416,1417,1417,1418,1418,1419,1419,1420,1420,1421,1421,1422,1422,1423,1423,1424,1424,1425,1425,1426,1426,1427,1427,1428,1428,1429,1429,1430,1430,1431,1431,1432,1432,1433,1433,1434,1434,1435,1435,1436,1436,1437,1437,1438,1438,1439,1439,1440,1440,1441,1441,1442,1442,1443,1443,1444,1444,1445,1445,1446,1446,1447,1447,1448,1448,1449,1449,1450,1450,1451,1451,1452,1452,1453,1453,1454,1454,1455,1455,1456,1456,1457,1457,1458,1458,1459,1459,1460,1460,1461,1461,1462,1462,1463,1463,1464,1464,1465,1465,1466,1466,1467,1467,1468,1468,1469,1469,1470,1470,1471,1471,1472,1472,1473,1473,1474,1474,1475,1475,1476,1476,1477,1477,1478,1478,1479,1479,1480,1480,1481,1481,1482,1482,1483,1483,1484,1484,1485,1485,1486,1486,1487,1487,1488,1488,1489,1489,1490,1490,1491,1491,1492,1492,1493,1493,1494,1494,1495,1495,1496,1496,1497,1497,1498,1498,1499,1499,1500,1500,1501,1501,1502,1502,1503,1503,1504,1504,1505,1505,1506,1506,1507,1507,1508,1508,1509,1509,1510,1510,1511,1511,1512,1512,1513,1513,1514,1514,1831,1831,1832,1832,1833,1833,1834,1834,1835,1835,1836,1836,1837,1837,1838,1838,1839,1839,1840,1840,1841,1841,1842,1842,1843,1843,1844,1844,1845,1845,1846,1846,1847,1847,1848,1848,1849,1849,1850,1850,1851,1851,1852,1852,1853,1853,1854,1854,1855,1855,1856,1856,1857,1857,1858,1858,1859,1859,1860,1860,1861,1861,1862,1862,1863,1863,1864,1864,1865,1865,1866,1866,1867,1867,1868,1868,1869,1869,1870,1870,1871,1871,1872,1872,1873,1873,1874,1874,1875,1875,1876,1876,1877,1877,1878,1878,1879,1879,1880,1880,1881,1881,1882,1882,1883,1883,1884,1884,1885,1885,1886,1886,1887,1887,1888,1888,1889,1889,1890,1890,1891,1891,1892,1892,1893,1893,1894,1894,1895,1895,1896,1896,1897,1897,1898,1898,1899,1899,1900,1900,1901,1901,1902,1902,1903,1903,1904,1904,1905,1905,1906,1906,1907,1907,1908,1908,1909,1909,1910,1910,1911,1911,1912,1912,1913,1913,1914,1914,1915,1915,1916,1916,1917,1917,1918,1918,1919,1919,1920,1920,1921,1921,1922,1922,1923,1923,1924,1924,1925,1925,1926,1926,1927,1927,1928,1928,1929,1929,1930,1930,1931,1931,1932,1932,1933,1933,1934,1934,1935,1935,1936,1936,1937,1937,1938,1938,1939,1939,1940,1940,1941,1941,1942,1942,1943,1943,1944,1944,1945,1945,1946,1946,1947,1947,1948,1948,1949,1949,1950,1950,1951,1951,1952,1952,1953,1953,1954,1954,1955,1955,1956,1956,1957,1957,1958,1958,1959,1959,1960,1960,1961,1961,1962,1962,1963,1963,1964,1964,1965,1965,1966,1966,1967,1967,1968,1968,1969,1969,1970,1970,1971,1971,1972,1972,1973,1973,1974,1974,1975,1975,1976,1976,1977,1977,1978,1978,1979,1979,1980,1980,1981,1981,1982,1982,1983,1983,1984,1984,1985,1985,1986,1986,1987,1987,1988,1988,1989,1989,1990,1990,1991,1991,1992,1992,1993,1993,1994,1994,1995,1995,1996,1996,1997,1997,1998,1998,1999,1999,2000,2000,2001,2001,2002,2002,2003,2003,2004,2004,2005,2005,2006,2006,2007,2007,2008,2008,2009,2009,2010,2010,2011,2011,2012,2012,2013,2013,2014,2014,2015,2015,2016,2016,2017,2017,2018,2018,2019,2019,2020,2020,2021,2021,2022,2022,2023,2023,2024,2024,2025,2025,2026,2026,2027,2027,2028,2028,2029,2029,2030,2030,2031,2031,2032,2032,2033,2033,2034,2034,2035,2035,2036,2036,2037,2037,2038,2038,2039,2039,2040,2040,2041,2041,2042,2042,2043,2043,2044,2044,2045,2045,2046,2046,2047,2047,2048,2048,2049,2049,2050,2050,2051,2051,2052,2052,2053,2053,2054,2054,2055,2055,2056,2056,2057,2057,2058,2058,2059,2059,2060,2060,2061,2061,2062,2062,2063,2063,2064,2064,2065,2065,2066,2066,2067,2067,2068,2068,2069,2069,2070,2070,2071,2071,2072,2072,2073,2073,2074,2074,2075,2075,2076,2076,2077,2077,2078,2078,2079,2079,2080,2080,2081,2081,2082,2082,2083,2083,2084,2084,2085,2085,2086,2086,2087,2087,2088,2088,2089,2089,2090,2090,2091,2091,2092,2092,2093,2093,2094,2094,2095,2095,2096,2096,2097,2097,2098,2098,2099,2099,2100,2100,2101,2101,2102,2102,2103,2103,2104,2104,2105,2105,2106,2106,2107,2107,2108,2108,2109,2109,2110,2110,2111,2111,2112,2112,2113,2113,2114,2114,2115,2115,2116,2116,2117,2117,2118,2118,2119,2119,2120,2120,2121,2121,2122,2122,2123,2123,2124,2124,2125,2125,2126,2126,2127,2127,2128,2128,2129,2129,2130,2130,2131,2131,2132,2132,2133,2133,2134,2134,2135,2135,2136,2136,2137,2137,2138,2138,2139,2139,2140,2140,2141,2141,2142,2142,2143,2143,2144,2144,2145,2145,2146,2146,2147,2147,2148,2148,2149,2149,2150,2150,2151,2151,2152,2152,2153,2153,2154,2154,2155,2155,2156,2156,2157,2157,2158,2158,2159,2159,2160,2160,2161,2161,2162,2162,2163,2163,2164,2164,2165,2165,2166,2166,2167,2167,2168,2168,2169,2169,2170,2170,2171,2171,2172,2172,2173,2173,2174,2174,2175,2175,2176,2176,2177,2177,2178,2178,2179,2179,2180,2180,2181,2181,2182,2182,2183,2183,2184,2184,2185,2185,2186,2186,2187,2187,2188,2188,2189,2189,2190,2190,2191,2191,2192,2192,2193,2193,2194,2194,2195,2195,2196,2196,2197,2197,2198,2198,2495,2495,2496,2496,2497,2497,2498,2498,2499,2499,2500,2500,2501,2501,2502,2502,2503,2503,2504,2504,2505,2505,2506,2506,2507,2507,2508,2508,2509,2509,2510,2510,2511,2511,2512,2512,2513,2513,2514,2514,2515,2515,2516,2516,2517,2517,2518,2518,2519,2519,2520,2520,2521,2521,2522,2522,2523,2523,2524,2524,2525,2525,2526,2526,2527,2527,2528,2528,2529,2529,2530,2530,2531,2531,2532,2532,2533,2533,2534,2534,2535,2535,2536,2536,2537,2537,2538,2538,2539,2539,2540,2540,2541,2541,2542,2542,2543,2543,2544,2544,2545,2545,2546,2546,2547,2547,2548,2548,2549,2549,2550,2550,2551,2551,2552,2552,2553,2553,2554,2554,2555,2555,2556,2556,2557,2557,2558,2558,2559,2559,2560,2560,2561,2561,2562,2562,2563,2563,2564,2564,2565,2565,2566,2566,2567,2567,2568,2568,2569,2569,2570,2570,2571,2571,2572,2572,2573,2573,2574,2574,2575,2575,2576,2576,2577,2577,2578,2578,2579,2579,2580,2580,2581,2581,2582,2582,2583,2583,2584,2584,2585,2585,2586,2586,2587,2587,2588,2588,2589,2589,2590,2590,2591,2591,2592,2592,2593,2593,2594,2594,2595,2595,2596,2596,2597,2597,2598,2598,2599,2599,2600,2600,2601,2601,2602,2602,2603,2603,2604,2604,2605,2605,2606,2606,2607,2607,2608,2608,2609,2609,2610,2610,2611,2611,2612,2612,2613,2613,2614,2614,2615,2615,2616,2616,2617,2617,2618,2618,2619,2619,2620,2620,2621,2621,2622,2622,2623,2623,2624,2624,2625,2625,2626,2626,2627,2627,2628,2628,2629,2629,2630,2630,2631,2631,2632,2632,2633,2633,2634,2634,2635,2635,2636,2636,2637,2637,2638,2638,2639,2639,2640,2640,2641,2641,2642,2642,2643,2643,2644,2644,2645,2645,2646,2646,2647,2647,2648,2648,2649,2649,2650,2650,2651,2651,2652,2652,2653,2653,2654,2654,2655,2655,2656,2656,2657,2657,2658,2658,2659,2659,2660,2660,2661,2661,2662,2662,2663,2663,2664,2664,2665,2665,2666,2666,2667,2667,2668,2668,2669,2669,2670,2670,2671,2671,2672,2672,2673,2673,2674,2674,2675,2675,2676,2676,2677,2677,2678,2678,2679,2679,2680,2680,2681,2681,2682,2682,2683,2683,2684,2684,2685,2685,2686,2686,2687,2687,2688,2688,2689,2689,2690,2690,2691,2691,2692,2692,2693,2693,2694,2694,2695,2695,2696,2696,2697,2697,2698,2698,2699,2699,2700,2700,2701,2701,2702,2702,2703,2703,2704,2704,2705,2705,2706,2706,2707,2707,2708,2708,2709,2709,2710,2710,2711,2711,2712,2712,2713,2713,2714,2714,2715,2715,2716,2716,2717,2717,2718,2718,2719,2719,2720,2720,2721,2721,2722,2722,2723,2723,2724,2724,2725,2725,2726,2726,2727,2727,2728,2728,2729,2729,2730,2730,2731,2731,2732,2732,2733,2733,2734,2734,2735,2735,2736,2736,2737,2737,2738,2738,2739,2739,2740,2740,2741,2741,2742,2742,2743,2743,2744,2744,2745,2745,2746,2746,2747,2747,2748,2748,2749,2749,2750,2750,2751,2751,2752,2752,2753,2753,2754,2754,2755,2755,2756,2756,2757,2757,2758,2758,2759,2759,2760,2760,2761,2761,2762,2762,2763,2763,2764,2764,2765,2765,2766,2766,3231,3231,3232,3232,3233,3233,3234,3234,3235,3235,3236,3236,3237,3237,3238,3238,3239,3239,3240,3240,3241,3241,3242,3242,3243,3243,3244,3244,3245,3245,3246,3246,3247,3247,3248,3248,3249,3249,3250,3250,3251,3251,3252,3252,3253,3253,3254,3254,3255,3255,3256,3256,3257,3257,3258,3258,3259,3259,3260,3260,3261,3261,3262,3262,3263,3263,3264,3264,3265,3265,3266,3266,3267,3267,3268,3268,3269,3269,3270,3270,3271,3271,3272,3272,3273,3273,3274,3274,3275,3275,3276,3276,3277,3277,3278,3278,3279,3279,3280,3280,3281,3281,3282,3282,3283,3283,3284,3284,3285,3285,3286,3286,3287,3287,3288,3288,3289,3289,3290,3290,3291,3291,3292,3292,3293,3293,3294,3294,3295,3295,3296,3296,3297,3297,3298,3298,3299,3299,3300,3300,3301,3301,3302,3302,3303,3303,3304,3304,3305,3305,3306,3306,3307,3307,3308,3308,3309,3309,3310,3310,3311,3311,3312,3312,3313,3313,3314,3314,3315,3315,3316,3316,3317,3317,3318,3318,3319,3319,3320,3320,3321,3321,3322,3322,3323,3323,3324,3324,3325,3325,3326,3326,3327,3327,3328,3328,3329,3329,3330,3330,3331,3331,3332,3332,3333,3333,3334,3334,3335,3335,3336,3336,3337,3337,3338,3338,3339,3339,3340,3340,3341,3341,3342,3342,3343,3343,3344,3344,3345,3345,3346,3346,3347,3347,3348,3348,3349,3349,3350,3350,3351,3351,3352,3352,3353,3353,3354,3354,3355,3355,3356,3356,3357,3357,3358,3358,3359,3359,3360,3360,3361,3361,3362,3362,3363,3363,3364,3364,3365,3365,3366,3366,3367,3367,3368,3368,3369,3369,3370,3370,3371,3371,3372,3372,3373,3373,3374,3374,3375,3375,3376,3376,3377,3377,3378,3378,3379,3379,3380,3380,3381,3381,3382,3382,3383,3383,3384,3384,3385,3385,3386,3386,3387,3387,3388,3388,3389,3389,3390,3390);
 constant depth : intArray(nNodes-1 downto 0)  :=  (0,1,1,2,2,2,2,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11);
 constant iLeaf : intArray(nLeaves-1 downto 0)  :=  (591,592,593,594,595,596,597,598,599,600,601,602,603,604,605,606,607,608,609,610,611,612,613,614,615,616,617,618,619,620,621,622,623,624,625,626,627,628,629,630,631,632,633,634,635,636,637,638,639,640,641,642,643,644,645,646,647,648,649,650,651,652,653,654,655,656,657,658,659,660,661,662,663,664,665,666,667,668,669,670,671,672,673,674,675,676,677,678,679,680,681,682,683,684,685,686,687,688,689,690,691,692,693,694,695,696,697,698,699,700,701,702,703,704,705,706,707,708,709,710,711,712,713,714,715,716,717,718,719,720,721,722,723,724,725,726,727,728,729,730,731,732,1057,1058,1059,1060,1061,1062,1063,1064,1065,1066,1067,1068,1069,1070,1071,1072,1073,1074,1075,1076,1077,1078,1079,1080,1081,1082,1083,1084,1085,1086,1087,1088,1089,1090,1091,1092,1093,1094,1095,1096,1097,1098,1099,1100,1101,1102,1103,1104,1105,1106,1107,1108,1109,1110,1111,1112,1113,1114,1115,1116,1117,1118,1119,1120,1121,1122,1123,1124,1125,1126,1127,1128,1129,1130,1131,1132,1133,1134,1135,1136,1137,1138,1139,1140,1141,1142,1143,1144,1145,1146,1147,1148,1149,1150,1151,1152,1153,1154,1155,1156,1157,1158,1159,1160,1161,1162,1163,1164,1165,1166,1167,1168,1169,1170,1171,1172,1173,1174,1175,1176,1177,1178,1179,1180,1181,1182,1515,1516,1517,1518,1519,1520,1521,1522,1523,1524,1525,1526,1527,1528,1529,1530,1531,1532,1533,1534,1535,1536,1537,1538,1539,1540,1541,1542,1543,1544,1545,1546,1547,1548,1549,1550,1551,1552,1553,1554,1555,1556,1557,1558,1559,1560,1561,1562,1563,1564,1565,1566,1567,1568,1569,1570,1571,1572,1573,1574,1575,1576,1577,1578,1579,1580,1581,1582,1583,1584,1585,1586,1587,1588,1589,1590,1591,1592,1593,1594,1595,1596,1597,1598,1599,1600,1601,1602,1603,1604,1605,1606,1607,1608,1609,1610,1611,1612,1613,1614,1615,1616,1617,1618,1619,1620,1621,1622,1623,1624,1625,1626,1627,1628,1629,1630,1631,1632,1633,1634,1635,1636,1637,1638,1639,1640,1641,1642,1643,1644,1645,1646,1647,1648,1649,1650,1651,1652,1653,1654,1655,1656,1657,1658,1659,1660,1661,1662,1663,1664,1665,1666,1667,1668,1669,1670,1671,1672,1673,1674,1675,1676,1677,1678,1679,1680,1681,1682,1683,1684,1685,1686,1687,1688,1689,1690,1691,1692,1693,1694,1695,1696,1697,1698,1699,1700,1701,1702,1703,1704,1705,1706,1707,1708,1709,1710,1711,1712,1713,1714,1715,1716,1717,1718,1719,1720,1721,1722,1723,1724,1725,1726,1727,1728,1729,1730,1731,1732,1733,1734,1735,1736,1737,1738,1739,1740,1741,1742,1743,1744,1745,1746,1747,1748,1749,1750,1751,1752,1753,1754,1755,1756,1757,1758,1759,1760,1761,1762,1763,1764,1765,1766,1767,1768,1769,1770,1771,1772,1773,1774,1775,1776,1777,1778,1779,1780,1781,1782,1783,1784,1785,1786,1787,1788,1789,1790,1791,1792,1793,1794,1795,1796,1797,1798,1799,1800,1801,1802,1803,1804,1805,1806,1807,1808,1809,1810,1811,1812,1813,1814,1815,1816,1817,1818,1819,1820,1821,1822,1823,1824,1825,1826,1827,1828,1829,1830,2199,2200,2201,2202,2203,2204,2205,2206,2207,2208,2209,2210,2211,2212,2213,2214,2215,2216,2217,2218,2219,2220,2221,2222,2223,2224,2225,2226,2227,2228,2229,2230,2231,2232,2233,2234,2235,2236,2237,2238,2239,2240,2241,2242,2243,2244,2245,2246,2247,2248,2249,2250,2251,2252,2253,2254,2255,2256,2257,2258,2259,2260,2261,2262,2263,2264,2265,2266,2267,2268,2269,2270,2271,2272,2273,2274,2275,2276,2277,2278,2279,2280,2281,2282,2283,2284,2285,2286,2287,2288,2289,2290,2291,2292,2293,2294,2295,2296,2297,2298,2299,2300,2301,2302,2303,2304,2305,2306,2307,2308,2309,2310,2311,2312,2313,2314,2315,2316,2317,2318,2319,2320,2321,2322,2323,2324,2325,2326,2327,2328,2329,2330,2331,2332,2333,2334,2335,2336,2337,2338,2339,2340,2341,2342,2343,2344,2345,2346,2347,2348,2349,2350,2351,2352,2353,2354,2355,2356,2357,2358,2359,2360,2361,2362,2363,2364,2365,2366,2367,2368,2369,2370,2371,2372,2373,2374,2375,2376,2377,2378,2379,2380,2381,2382,2383,2384,2385,2386,2387,2388,2389,2390,2391,2392,2393,2394,2395,2396,2397,2398,2399,2400,2401,2402,2403,2404,2405,2406,2407,2408,2409,2410,2411,2412,2413,2414,2415,2416,2417,2418,2419,2420,2421,2422,2423,2424,2425,2426,2427,2428,2429,2430,2431,2432,2433,2434,2435,2436,2437,2438,2439,2440,2441,2442,2443,2444,2445,2446,2447,2448,2449,2450,2451,2452,2453,2454,2455,2456,2457,2458,2459,2460,2461,2462,2463,2464,2465,2466,2467,2468,2469,2470,2471,2472,2473,2474,2475,2476,2477,2478,2479,2480,2481,2482,2483,2484,2485,2486,2487,2488,2489,2490,2491,2492,2493,2494,2767,2768,2769,2770,2771,2772,2773,2774,2775,2776,2777,2778,2779,2780,2781,2782,2783,2784,2785,2786,2787,2788,2789,2790,2791,2792,2793,2794,2795,2796,2797,2798,2799,2800,2801,2802,2803,2804,2805,2806,2807,2808,2809,2810,2811,2812,2813,2814,2815,2816,2817,2818,2819,2820,2821,2822,2823,2824,2825,2826,2827,2828,2829,2830,2831,2832,2833,2834,2835,2836,2837,2838,2839,2840,2841,2842,2843,2844,2845,2846,2847,2848,2849,2850,2851,2852,2853,2854,2855,2856,2857,2858,2859,2860,2861,2862,2863,2864,2865,2866,2867,2868,2869,2870,2871,2872,2873,2874,2875,2876,2877,2878,2879,2880,2881,2882,2883,2884,2885,2886,2887,2888,2889,2890,2891,2892,2893,2894,2895,2896,2897,2898,2899,2900,2901,2902,2903,2904,2905,2906,2907,2908,2909,2910,2911,2912,2913,2914,2915,2916,2917,2918,2919,2920,2921,2922,2923,2924,2925,2926,2927,2928,2929,2930,2931,2932,2933,2934,2935,2936,2937,2938,2939,2940,2941,2942,2943,2944,2945,2946,2947,2948,2949,2950,2951,2952,2953,2954,2955,2956,2957,2958,2959,2960,2961,2962,2963,2964,2965,2966,2967,2968,2969,2970,2971,2972,2973,2974,2975,2976,2977,2978,2979,2980,2981,2982,2983,2984,2985,2986,2987,2988,2989,2990,2991,2992,2993,2994,2995,2996,2997,2998,2999,3000,3001,3002,3003,3004,3005,3006,3007,3008,3009,3010,3011,3012,3013,3014,3015,3016,3017,3018,3019,3020,3021,3022,3023,3024,3025,3026,3027,3028,3029,3030,3031,3032,3033,3034,3035,3036,3037,3038,3039,3040,3041,3042,3043,3044,3045,3046,3047,3048,3049,3050,3051,3052,3053,3054,3055,3056,3057,3058,3059,3060,3061,3062,3063,3064,3065,3066,3067,3068,3069,3070,3071,3072,3073,3074,3075,3076,3077,3078,3079,3080,3081,3082,3083,3084,3085,3086,3087,3088,3089,3090,3091,3092,3093,3094,3095,3096,3097,3098,3099,3100,3101,3102,3103,3104,3105,3106,3107,3108,3109,3110,3111,3112,3113,3114,3115,3116,3117,3118,3119,3120,3121,3122,3123,3124,3125,3126,3127,3128,3129,3130,3131,3132,3133,3134,3135,3136,3137,3138,3139,3140,3141,3142,3143,3144,3145,3146,3147,3148,3149,3150,3151,3152,3153,3154,3155,3156,3157,3158,3159,3160,3161,3162,3163,3164,3165,3166,3167,3168,3169,3170,3171,3172,3173,3174,3175,3176,3177,3178,3179,3180,3181,3182,3183,3184,3185,3186,3187,3188,3189,3190,3191,3192,3193,3194,3195,3196,3197,3198,3199,3200,3201,3202,3203,3204,3205,3206,3207,3208,3209,3210,3211,3212,3213,3214,3215,3216,3217,3218,3219,3220,3221,3222,3223,3224,3225,3226,3227,3228,3229,3230,3391,3392,3393,3394,3395,3396,3397,3398,3399,3400,3401,3402,3403,3404,3405,3406,3407,3408,3409,3410,3411,3412,3413,3414,3415,3416,3417,3418,3419,3420,3421,3422,3423,3424,3425,3426,3427,3428,3429,3430,3431,3432,3433,3434,3435,3436,3437,3438,3439,3440,3441,3442,3443,3444,3445,3446,3447,3448,3449,3450,3451,3452,3453,3454,3455,3456,3457,3458,3459,3460,3461,3462,3463,3464,3465,3466,3467,3468,3469,3470,3471,3472,3473,3474,3475,3476,3477,3478,3479,3480,3481,3482,3483,3484,3485,3486,3487,3488,3489,3490,3491,3492,3493,3494,3495,3496,3497,3498,3499,3500,3501,3502,3503,3504,3505,3506,3507,3508,3509,3510,3511,3512,3513,3514,3515,3516,3517,3518,3519,3520,3521,3522,3523,3524,3525,3526,3527,3528,3529,3530,3531,3532,3533,3534,3535,3536,3537,3538,3539,3540,3541,3542,3543,3544,3545,3546,3547,3548,3549,3550,3551,3552,3553,3554,3555,3556,3557,3558,3559,3560,3561,3562,3563,3564,3565,3566,3567,3568,3569,3570,3571,3572,3573,3574,3575,3576,3577,3578,3579,3580,3581,3582,3583,3584,3585,3586,3587,3588,3589,3590,3591,3592,3593,3594,3595,3596,3597,3598,3599,3600,3601,3602,3603,3604,3605,3606,3607,3608,3609,3610,3611,3612,3613,3614,3615,3616,3617,3618,3619,3620,3621,3622,3623,3624,3625,3626,3627,3628,3629,3630,3631,3632,3633,3634,3635,3636,3637,3638,3639,3640,3641,3642,3643,3644,3645,3646,3647,3648,3649,3650,3651,3652,3653,3654,3655,3656,3657,3658,3659,3660,3661,3662,3663,3664,3665,3666,3667,3668,3669,3670,3671,3672,3673,3674,3675,3676,3677,3678,3679,3680,3681,3682,3683,3684,3685,3686,3687,3688,3689,3690,3691,3692,3693,3694,3695,3696,3697,3698,3699,3700,3701,3702,3703,3704,3705,3706,3707,3708,3709,3710,3711,3712,3713,3714,3715,3716,3717,3718,3719,3720,3721,3722,3723,3724,3725,3726,3727,3728,3729,3730,3731,3732,3733,3734,3735,3736,3737,3738,3739,3740,3741,3742,3743,3744,3745,3746,3747,3748,3749,3750,3751,3752,3753,3754,3755,3756,3757,3758,3759,3760,3761,3762,3763,3764,3765,3766,3767,3768,3769,3770,3771,3772,3773,3774,3775,3776,3777,3778,3779,3780,3781,3782,3783,3784,3785,3786,3787,3788,3789,3790,3791,3792,3793,3794,3795,3796,3797,3798,3799,3800,3801,3802,3803,3804,3805,3806,3807,3808,3809,3810,3811,3812,3813,3814,3815,3816,3817,3818,3819,3820,3821,3822,3823,3824,3825,3826,3827,3828,3829,3830,3831,3832,3833,3834,3835,3836,3837,3838,3839,3840,3841,3842,3843,3844,3845,3846,3847,3848,3849,3850,3851,3852,3853,3854,3855,3856,3857,3858,3859,3860,3861,3862,3863,3864,3865,3866,3867,3868,3869,3870,3871,3872,3873,3874,3875,3876,3877,3878,3879,3880,3881,3882,3883,3884,3885,3886,3887,3888,3889,3890,3891,3892,3893,3894,3895,3896,3897,3898,3899,3900,3901,3902,3903,3904,3905,3906,3907,3908,3909,3910,3911,3912,3913,3914,3915,3916,3917,3918,3919,3920,3921,3922,3923,3924,3925,3926,3927,3928,3929,3930,3931,3932,3933,3934,3935,3936,3937,3938,3939,3940,3941,3942,3943,3944,3945,3946,3947,3948,3949,3950,3951,3952,3953,3954,3955,3956,3957,3958,3959,3960,3961,3962,3963,3964,3965,3966,3967,3968,3969,3970,3971,3972,3973,3974,3975,3976,3977,3978,3979,3980,3981,3982,3983,3984,3985,3986,3987,3988,3989,3990,3991,3992,3993,3994,3995,3996,3997,3998,3999,4000,4001,4002,4003,4004,4005,4006,4007,4008,4009,4010,4011,4012,4013,4014,4015,4016,4017,4018,4019,4020,4021,4022,4023,4024,4025,4026,4027,4028,4029,4030,4031,4032,4033,4034,4035,4036,4037,4038,4039,4040,4041,4042,4043,4044,4045,4046,4047,4048,4049,4050,4051,4052,4053,4054,4055,4056,4057,4058,4059,4060,4061,4062,4063,4064,4065,4066,4067,4068,4069,4070,4071,4072,4073,4074,4075,4076,4077,4078,4079,4080,4081,4082,4083,4084,4085,4086,4087,4088,4089,4090,4091,4092,4093,4094);
constant value     : tyArray(nNodes-1 downto 0) := to_tyArray(value_int);
constant threshold  : txArray(nNodes-1 downto 0) := to_txArray(threshold_int);
 end Arrays0_0000;
